`define DELAY 20
module alu_32bit_testbench();

reg [31:0] a, b;
reg [2:0] op_code;
wire [31:0] result;
wire c_out, Z;

alu_32bit test_alu_33bit (a, b, op_code, result, c_out, Z);

initial begin
	///////////////////////////////////AND
	a=32'b11110000111100001111111100000000;
	b=32'b11111111000011110000111100000000;
	op_code=3'b000;
	#`DELAY;
	
	///////////////////////////////////OR
	a=32'b11110000111100001111111100000000;
	b=32'b11111111000011110000111100000000;
	op_code=3'b001;
	#`DELAY;
	
	///////////////////////////////////ADD
	a=32'b00000000000000001111111100000000;
	b=32'b00000000000011110000111100000000;
	op_code=3'b010;
	#`DELAY;
	
	a=32'b10001111111110001111111100000000;
	b=32'b10111111110011110000111100111100;
	op_code=3'b010;
	#`DELAY;
	
	a=32'b00000000111100001111111100000000;
	b=32'b11111111000011110000111100000000;
	op_code=3'b010;
	#`DELAY;
	
	///////////////////////////////////SUBTRACT
	a=32'b00000000000000001111111100000000;
	b=32'b00000000000011110000111100000000;
	op_code=3'b110;
	#`DELAY;
	
	a=32'b00001010010100001111111100000000;
	b=32'b00000000000011110000111100000000;
	op_code=3'b110;
	#`DELAY;
	
	a=32'b11111000000000000000000000000000;
	b=32'b10000111100000000000000000000000;
	op_code=3'b110;
	#`DELAY;
	
	a=32'b10000111100000000000000000000000;
	b=32'b11111000000000000000000000000000;
	op_code=3'b110;
	#`DELAY;
	
	a=32'b11111000011110000011110000000000;
	b=32'b00011000000110000011110000000000;
	op_code=3'b110;
	#`DELAY;
	
	a=32'b00000000011100001000011110000000;
	b=32'b11111000011110000000111100011110;
	op_code=3'b110;
	#`DELAY;
	
	///////////////////////////////////XOR
	a=32'b11110000111100001111111100000000;
	b=32'b11111111000011110000111100000000;
	op_code=3'b011;
	#`DELAY;
	
	////////////////////////////////////Zero Bit
	a=32'b11110000111100001111111100000000;
	b=32'b11111111000011110000111100000000;
	op_code=3'b110;
	#`DELAY;
	
	a=32'b00000000000000000000000000000000;
	b=32'b00000000000000000000000000000000;
	op_code=3'b110;
	#`DELAY;
	
	a=32'b11111111111111111111111111111111;
	b=32'b11111111111111111111111111111111;
	op_code=3'b110;
	#`DELAY;
	
	
end

initial begin
	$monitor("a=%32b, b=%32b, op_code=%3b, result=%32b, c_out=%1b, Z=%1b ",a, b, op_code, result, c_out, Z);
end


endmodule

/*
ALUop		Function
000		AND
001		OR
010		ADD
110		SUBTRACT
011		XOR
*/
